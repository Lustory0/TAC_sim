** Profile: "SCHEMATIC1-sim_psp"  [ c:\cds_spb_home\cdssetup\project4\project4-pspicefiles\schematic1\sim_psp.sim ] 

** Creating circuit file "sim_psp.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2.65u 2.35u 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.OPTIONS ABSTOL= 1.0n
.OPTIONS ITL4= 1000
.OPTIONS RELTOL= 0.01
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
